library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fir_coeffs_pkg is
	-- Jednostavan tip za niz real koeficijenata (dužina se zadaje pri deklaraciji konstante)
	type real_vec_t is array (natural range <>) of real;

	------------------------------------------------------------------------------
	-- STAGE 0 (N = 42)  — tvoji postojeći koeficijenti
	------------------------------------------------------------------------------
	constant FIR0_N : natural := 42;

	constant FIR0_PH0_R : real_vec_t(0 to FIR0_N-1) := (
		0.000014291322,
		-0.000039516421,
		0.000091072642,
		-0.000183517720,
		0.000337020847,
		-0.000578304995,
		0.000940386412,
		-0.001464323420,
		0.002199199950,
		-0.003204611510,
		0.004552420300,
		-0.006332841260,
		0.008663313130,
		-0.011708605900,
		0.015718495800,
		-0.021111531700,
		0.028669391700,
		-0.040069744000,
		0.059694815000,
		-0.103678482000,
		0.317492818000,
		0.317492818000,
		-0.103678482000,
		0.059694815000,
		-0.040069744000,
		0.028669391700,
		-0.021111531700,
		0.015718495800,
		-0.011708605900,
		0.008663313130,
		-0.006332841260,
		0.004552420300,
		-0.003204611510,
		0.002199199950,
		-0.001464323420,
		0.000940386412,
		-0.000578304995,
		0.000337020847,
		-0.000183517720,
		0.000091072642,
		-0.000039516421,
		0.000014291322
	);

	constant FIR0_PH1_R : real_vec_t(0 to FIR0_N-1) := (
		0.000000000000,
		-0.000000125470,
		0.000000200697,
		-0.000000503721,
		0.000000828311,
		-0.000001458836,
		0.000002191536,
		-0.000003306305,
		0.000004591620,
		-0.000006307723,
		0.000008197802,
		-0.000010484277,
		0.000012878196,
		-0.000015551202,
		0.000018184220,
		-0.000020897352,
		0.000023348090,
		-0.000025659990,
		0.000027483840,
		-0.000028956372,
		0.000029782526,
		0.499967636000,
		0.000029782526,
		-0.000028956372,
		0.000027483840,
		-0.000025659990,
		0.000023348090,
		-0.000020897352,
		0.000018184220,
		-0.000015551202,
		0.000012878196,
		-0.000010484277,
		0.000008197802,
		-0.000006307723,
		0.000004591620,
		-0.000003306305,
		0.000002191536,
		-0.000001458836,
		0.000000828311,
		-0.000000503721,
		0.000000200697,
		-0.000000125470
	);

	------------------------------------------------------------------------------
	-- STAGE 1 — koeficijenti iz tvojih fajlova (ph0: 10 tapova, ph1: 9 tapova)
	------------------------------------------------------------------------------
	constant FIR1_N : natural := 10;

	constant FIR1_PH0_R : real_vec_t(0 to FIR1_N-1) := (
		0.000745880558,
		-0.005654152930,
		0.023419375400,
		-0.074944555800,
		0.306435005000,
		0.306435005000,
		-0.074944555800,
		0.023419375400,
		-0.005654152930,
		0.000745880558
	);

	constant FIR1_PH1_R : real_vec_t(0 to FIR1_N-1) := (
		0.000000000000,
		-0.000000000000,
		0.000000000000,
		-0.000000000000,
		0.499996896000,
		-0.000000000000,
		0.000000000000,
		-0.000000000000,
		0.000000000000,
		0.0
	);

	------------------------------------------------------------------------------
	-- STAGE 2 — koeficijenti iz tvojih fajlova (ph0: 6 tapova, ph1: 5 tapova)
	------------------------------------------------------------------------------
	constant FIR2_N : natural := 6;

	constant FIR2_PH0_R : real_vec_t(0 to FIR2_N-1) := (
		0.006730474570,
		-0.051299722400,
		0.294570558000,
		0.294570558000,
		-0.051299722400,
		0.006730474570
	);

	constant FIR2_PH1_R : real_vec_t(0 to FIR2_N-1) := (
		0.000018084556,
		-0.000062439061,
		0.500086089000,
		-0.000062439061,
		0.000018084556,
		0.0
	);

end package fir_coeffs_pkg;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package lut_pkg is
	-- VHDL-2008: unconstrained row; svaka tabela ima svoj N (broj kolona)
	subtype row_t is std_logic_vector;              -- (N-1 downto 0)
	type    rom16_t is array (0 to 15) of row_t;    -- 16 nivoa: +7 .. -8

	--------------------------------------------------------------------
	-- LUT1  (preuzeto iz LUT1.txt, izbačen prvi red = +8)
	-- 16 vrsta: +7 .. -8 ; N = 16 kolona
	--------------------------------------------------------------------
	constant LUT1_ROM : rom16_t := (
		0	=> "0111111111111111",
		1	=> "0111111111111101",
		2	=> "0101111111111101",
		3	=> "0101111111110101",
		4	=> "0101111111101010",
		5	=> "0101011111010101",
		6	=> "0101011101010101",
		7	=> "0101010101010101",
		8	=> "0101010001010101",
		9	=> "0101000001010101",
		10	=> "0101000000010101",
		11	=> "0101000000000101",
		12	=> "0100000000000101",
		13	=> "0100000000000001",
		14	=> "0000000000000001",
		15	=> "0000000000000000"
	);
	constant LUT1_LEN : natural := 16;	-- kolona

	--------------------------------------------------------------------
	-- LUT2  (preuzeto iz LUT2.txt, izbačen prvi red = +8)
	-- 16 vrsta: +7 .. -8 ; N = 32 kolone
	--------------------------------------------------------------------
	constant LUT2_ROM : rom16_t := (
		0	=> "01111111111111111111111111111110",
		1	=> "01111111111111011011111111111110",
		2	=> "01011111111111011011111111111010",
		3	=> "01011111111101011010111111111010",
		4	=> "01011111110101011010101111111010",
		5	=> "01010111110101011010101111101010",
		6	=> "01010111010101011010101011101010",
		7	=> "01010101010101011010101010101010",
		8	=> "10101000101010100101010100010101",
		9	=> "10101000001010100101010000010101",
		10	=> "10100000001010100101010000000101",
		11	=> "10100000000010100101000000000101",
		12	=> "10100000000000100100000000000101",
		13	=> "10000000000000100100000000000001",
		14	=> "10000000000000000000000000000001",
		15	=> "00000000000000000000000000000000"
	);
	constant LUT2_LEN : natural := 32;	-- kolona

	--------------------------------------------------------------------
	-- LUT3  (preuzeto iz LUT3.txt, izbačen prvi red = +8)
	-- 16 vrsta: +7 .. -8 ; N = 32 kolone
	--------------------------------------------------------------------
	constant LUT3_ROM : rom16_t := (
		0	=> "11111101111111111111111110111111",
		1	=> "11101111111101111110111111110111",
		2	=> "11101111001111111111110011110111",
		3	=> "10111110011111011011111001111101",
		4	=> "11110000111011111111011100001111",
		5	=> "10101101101101100110110110110101",
		6	=> "11100001010011111111001010000111",
		7	=> "01101001100101100110100110010110",
		8	=> "00011110101100000000110101111000",
		9	=> "01010010010010011001001001001010",
		10	=> "00001111000100000000100011110000",
		11	=> "01000001100000100100000110000010",
		12	=> "00010000110000000000001100001000",
		13	=> "00010000000010000001000000001000",
		14	=> "00000010000000000000000100000000",
		15	=> "00000000000000000000000000000000"
	);
	constant LUT3_LEN : natural := 32;	-- kolona

	--------------------------------------------------------------------
	-- LUT4  (mid-rise; preuzeto iz LUT4.txt)
	-- 16 vrsta: +7 .. -8 ; N = 15 kolona
	--------------------------------------------------------------------
	constant LUT4_ROM : rom16_t := (
		0	=> "111111111111111",
		1	=> "111111101111111",
		2	=> "111011111110111",
		3	=> "110111101111011",
		4	=> "101111010111101",
		5	=> "101101101101101",
		6	=> "101010111010101",
		7	=> "100110101011001",
		8	=> "011001010100110",
		9	=> "010101000101010",
		10	=> "010010010010010",
		11	=> "010000101000010",
		12	=> "001000010000100",
		13	=> "000100000001000",
		14	=> "000000010000000",
		15	=> "000000000000000"
	);
	constant LUT4_LEN : natural := 15;	-- kolona

	--------------------------------------------------------------------
	-- LUT5  (mid-rise; preuzeto iz LUT5.txt)
	-- 16 vrsta: +7 .. -8 ; N = 19 kolona
	--------------------------------------------------------------------
	constant LUT5_ROM : rom16_t := (
		0	=> "1111011111111101111",
		1	=> "1101111110111111011",
		2	=> "1110011111111100111",
		3	=> "1101011110111101011",
		4	=> "1011011101011101101",
		5	=> "1011001110111001101",
		6	=> "1010101011101010101",
		7	=> "0101111000001111010",
		8	=> "1010000111110000101",
		9	=> "0101010100010101010",
		10	=> "0100110001000110010",
		11	=> "0100100010100010010",
		12	=> "0010100001000010100",
		13	=> "0001100000000011000",
		14	=> "0010000001000000100",
		15	=> "0000100000000010000"
	);
	constant LUT5_LEN : natural := 19;	-- kolona
	
	--------------------------------------------------------------------
	-- API funkcije (deklaracije)
	--------------------------------------------------------------------
	function lut_len(id : integer) return natural;
	function get_row(id : integer; idx : integer) return row_t;
	
	-- mapiranje ulaza: [-2^(W-1) .. 2^(W-1)-1] -> 0..2^W-1 uz flip
	-- prima vektor proizvoljne širine i vraća unsigned iste širine
	function map_row_index(d : std_logic_vector) return unsigned;

end package;

package body lut_pkg is

  function lut_len(id : integer) return natural is
  begin
    case id is
      when 1      => return LUT1_LEN;
      when 2      => return LUT2_LEN;
      when 3      => return LUT3_LEN;
      when 4      => return LUT4_LEN;
      when 5      => return LUT5_LEN;
      when others => return LUT1_LEN;
    end case;
  end function;

  function get_row(id : integer; idx : integer) return row_t is
  begin
    case id is
      when 1      => return LUT1_ROM(idx);
      when 2      => return LUT2_ROM(idx);
      when 3      => return LUT3_ROM(idx);
      when 4      => return LUT4_ROM(idx);
      when 5      => return LUT5_ROM(idx);
      when others => return LUT1_ROM(idx);
    end case;
  end function;

  function map_row_index(d : std_logic_vector) return unsigned is
    constant W    : natural := d'length;
    constant BIAS : signed(d'range) := to_signed(2**(W-1), W);
    variable u    : unsigned(d'range);
  begin
    -- shift u 0..2^W-1
    u := unsigned(signed(d) + BIAS);
    -- flip: (2^W-1) - u  == bitwise not za tačnu širinu
    return not u;
  end function;

end package body;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package deltaSigma_pkg is

	constant C_X_UPPER	: integer	:= 3;
	constant C_X_LOWER	: integer	:= -8;
	constant C_Y_UPPER	: integer	:= 4;
	constant C_Y_LOWER	: integer	:= 0;
	

end package deltaSigma_pkg;